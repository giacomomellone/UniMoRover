----------------------------------------------------------------------------------
-- PSE 2016/2017
-- Students: Mazzocchi, Mellone, Pistoni, Truffellini, Vidoni

-- Module Name:    Display7 - Behavioral 
-- Description:    7 segment display showing LH, RH, UP or DOWN and HORN according
-- to pushed button
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Display7 is
    Port ( BTN : in  STD_LOGIC_VECTOR (4 downto 0);
           SEG : out  STD_LOGIC_VECTOR (7 downto 0);
			  AN : out  STD_LOGIC_VECTOR (3 downto 0);
			  CLK : in STD_LOGIC; -- 5 MHz clock, generated by PLL
			  COMMAND : out STD_LOGIC_VECTOR (7 downto 0) -- Byte sent to PIC18LF25K80
			 );
end Display7;

-- Font ROM
-- SEG <= "10001001"; -- H
-- SEG <= "10100001"; -- d
-- SEG <= "11000001"; -- U
-- SEG <= "10001100"; -- P
-- SEG <= "10100011"; -- o
-- SEG <= "11100011"; -- u/w
-- SEG <= "10101011"; -- n
-- SEG <= "11000111"; -- L
-- SEG <= "10101111"; -- r
-- SEG <= "10000110"; -- E
-- SEG <= "10000111"; -- t
-- SEG <= "10001110"; -- F
-- SEG <= "10111111"; -- -

architecture Behavioral of Display7 is

	signal cnt : Integer range 0 to 2147483640:= 0;
	-- This counter is needed to count the clock period for which one has to illuminate each
	-- anode in order to provide the human eye with the information.
	
begin

process(CLK)
begin
AN <= "1111";
if(CLK'event and CLK='1')then
	cnt <= cnt+1;
	
-- UP command
	if (BTN(0)='1' AND BTN(1)='0' AND BTN(2)='0' AND BTN(3)='0' AND BTN(4)='0') then
		COMMAND <= X"55"; -- ascii = U
		if cnt<10000 then
			AN <= "0111";
			SEG <= "11000001"; -- U
		elsif (cnt>=10000 AND cnt<20000) then
			AN <= "1011";
			SEG <= "10001100"; -- P
		else
			cnt <= 0;
		end if;
		
-- LEFT command
	elsif (BTN(0)='0' AND BTN(1)='1' AND BTN(2)='0' AND BTN(3)='0' AND BTN(4)='0') then
		COMMAND <= X"4C"; -- ascii = L
		if cnt<10000 then
			AN <= "0111";
			SEG <= "11000111"; -- L
		elsif (cnt>=10000 AND cnt<20000) then
			AN <= "1011";
			SEG <= "10000110"; -- E
		elsif (cnt>=20000 AND cnt<30000) then
			AN <= "1101";
			SEG <= "10001110"; -- F
		elsif (cnt>=30000 AND cnt<40000) then
			AN <= "1110";
			SEG <= "10000111"; -- t
		else
			cnt <= 0;
		end if;

-- RIGHT command
	elsif (BTN(0)='0' AND BTN(1)='0' AND BTN(2)='0' AND BTN(3)='1' AND BTN(4)='0') then
		COMMAND <= X"52"; -- ascii = R
		if cnt<10000 then
			AN <= "0111";
			SEG <= "10101111"; -- r
		elsif (cnt>=10000 AND cnt<20000) then
			AN <= "1011";
			SEG <= "10001001"; -- H
		else
			cnt <= 0;
		end if;

-- DOWN command
	elsif (BTN(0)='0' AND BTN(1)='0' AND BTN(2)='1' AND BTN(3)='0' AND BTN(4)='0') then
		COMMAND <= X"44"; -- ascii = D
		if cnt<10000 then
			AN <= "0111";
			SEG <= "10100001"; -- d
		elsif (cnt>=10000 AND cnt<20000) then
			AN <= "1011";
			SEG <= "10100011"; -- o
		elsif (cnt>=20000 AND cnt<30000) then
			AN <= "1101";
			SEG <= "11100011"; -- w
		elsif (cnt>=30000 AND cnt<40000) then
			AN <= "1110";
			SEG <= "10101011"; -- n
		else
			cnt <= 0;
		end if;

-- HORN command
	elsif (BTN(0)='0' AND BTN(1)='0' AND BTN(2)='0' AND BTN(3)='0' AND BTN(4)='1') then
		COMMAND <= X"48"; -- ascii = H
		if cnt<10000 then
			AN <= "0111";
			SEG <= "10001001"; -- H
		elsif (cnt>=10000 AND cnt<20000) then
			AN <= "1011";
			SEG <= "10100011"; -- o
		elsif (cnt>=20000 AND cnt<30000) then
			AN <= "1101";
			SEG <= "10101111"; -- r
		elsif (cnt>=30000 AND cnt<40000) then
			AN <= "1110";
			SEG <= "10101011"; -- n
		else
			cnt <= 0;
		end if;
		
		
-- UP-HORN command
-- It could be useful to have this command in case of humans in front of the vehicle
	elsif (BTN(0)='1' AND BTN(1)='0' AND BTN(2)='0' AND BTN(3)='0' AND BTN(4)='1') then
		COMMAND <= X"68"; -- ascii = h
		if cnt<10000 then
			AN <= "0111";
			SEG <= "11000001"; -- U
		elsif (cnt>=10000 AND cnt<20000) then
			AN <= "1011";
			SEG <= "10001100"; -- P
		elsif (cnt>=20000 AND cnt<30000) then
			AN <= "1101";
			SEG <= "10111111"; -- -
		elsif (cnt>=30000 AND cnt<40000) then
			AN <= "1110";
			SEG <= "10001001"; -- H
		else
			cnt <= 0;
		end if;
		
-- In all other cases, like pressing together 3 buttons and presing nothing
	-- STOP - S
	else
		COMMAND <= X"53"; -- ascii = S
		SEG <= "11111111";
		AN <= "1111";
	end if;
	-- STOP - S
	if (BTN(0)='0' AND BTN(1)='0' AND BTN(2)='0' AND BTN(3)='0' AND BTN(4)='0') then
		COMMAND <= X"53"; -- ascii = S
		SEG <= "11111111";
		AN <= "1111";
		cnt <= 0;
	end if;
end if;
end process;
end Behavioral;
